module Decoder3to8(x2, x1, x0, w0, w1, w2, w3, w4, w5, w6, w7, en);
	input x2, x1, x0, en;
	output reg w0, w1, w2, w3, w4, w5, w6, w7;
	
	always @(x2 or x1 or x0)
	begin
		case ({en, x2, x1, x0})
			4'b0000: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b0001: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b0010: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b0011: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b0100: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b0101: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b0110: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b0111: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000000;
			4'b1000: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000001;
			4'b1001: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000010;
			4'b1010: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00000100;
			4'b1011: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00001000;
			4'b1100: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00010000;
			4'b1101: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b00100000;
			4'b1110: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b01000000;
			4'b1111: {w7, w6, w5, w4, w3, w2, w1, w0} = 8'b10000000;
		endcase
	end
endmodule
